module konstanta (output c, input a);
   assign c = 1 | a;  
endmodule