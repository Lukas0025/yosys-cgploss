module xordecoder (input a,
                  output [127:0] out);
	assign out = {   a ^ a,
			 a ^ a ^ a,
			 a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a,
			 a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a ^ a};
endmodule