module empty_tb; 
  initial begin
  end
endmodule